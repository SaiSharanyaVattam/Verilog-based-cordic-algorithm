module testbench();
reg [31:0] zin;
wire [31:0]sinho, cosho, tanho;
cordic_sin_cos UUT(zin, sinho, cosho, tanho);
initial begin
zin=32'b01000000000000000000000000000000;
//zin=32'b00111111100000000000000000000000;//1
//zin=32'b10111111011001100110011001100110;//0.9
//zin=32'b00111111001100110011001100110011;//0.7
//zin=32'b01000000000000000000000000000000;//45
//zin=32'b01000010001101000000000000000000;//30
end
endmodule
